BZh91AY&SYcc �_�Py����߰����`���5X���:  dɓ��&	�F�!��&L��L �0L�0�M��L@ �     ���j4�ɠhb&#h��z�)&�A4������  ���L&�4��&A����&��ښy�P�i��U�@��Jp|��e
4�KO����#橢�� �B�Ԙ��%���e��.(Y!ZJOW��o�*lg'�O5L����f�K����Q$�=3��Ek8N�(�(/�d��&�s2��h��������k}�TÓ�n�&F%g87*R��KK�fŘJ��T��	gn��t�����DU��{����,���s�6�dT�*UUQ^w��lcoV�>��J4
df�1Fa	{,�_/3f�dúҿej���0�h^���^��Tw��b-4##;9�ʭ
11m��x[
K���*@aCK�� -���@�9�d�[R(���f�H�k��e���Z�4qDC�&�y�sw��$!B^IHI!�IwU���_J	�BB�)S2�P8�P�AF4��@$:H$��!j�(Ad3�'�H�A�J0�D(d�OX>T�6�=L�:M�����<
T*l�V�{x�+�L��3ׯ��qln{c�F�BV1�k�0�2�)��*�;�8��3��m���R�{�߯����*jd]��.�'6N���r��̗v�s~l���$��n}/r��r��d�bX�A
�D�U�����<�ys��a���rY0��q]�����\���b�����z��]e؛T]�;.FNH�k��%�"����<�ڥ�}�\F���e�v����:nnVl:p`�E��g��g����`���e&��ر%�ԓ�1bּ��c�fB���sQ��&2ȱXԪ���۽*h`��:d�d�E�eJn�̚ڤ�$�)�41���܋wܷvN�(�D]yd�]:���˔|��Ǳ1����SR\������W'q�������B��v'������ϵŋq�!�䢪(��?g$��I"�F����K�In3�EC��Z�9ҵ�*yT�����`3,��]�51�L'
��Y)�7�"�5�bT]�?� �2�ZlhR^)d���,�b��j�c5,��x�v	b�ף�Z4=�rE�C���B���AҎ��dS�[��I����)�{6��v��7�wL\6Λ,�c����P��%!�X{�s�w7TN-LU*B�s���ns�a]V���"�IG�b㑱�3t;��gcŋtq�h��7p*d��E�yz]s�	)]�N�X�_��,�Rlwg�l�f)��_s$k��Ŏ�����Š�e2�N�d3ll�&�/�J���M�4oT�]��^n����ٴkN�5��[F��r,6<X��p�����s0.�y�`�}�y�N�����;��'���J����:4���u)���א�*)F-m��H�
b�,`