BZh91AY&SY��#� �_�Py����������`� �4    jM=CF�hɠ4dh  �<C$ʞj� 4�4ɐ ���&L��L �0L�0�2d�b`ɂd ф``8ɓ&# &L �# C � @�0L��hѪ~��=��mO?E1��_��ILB \�?$�h�ͮ#b��"}������y\4�0APC�Ђ�4�i%V��d1hG��E�]ۄ~z������G�R��uׁR�>j>-I:C�L�t����;X� �d�̃M�IJr��4]��y���)�萘QY˘���ю2�����I��Tԧ:��I�u�Y�	�`x Y�g��.��$�{��Ep#G!ݠ;��Ik&M�M??�Ѫ�ذ�+Ĉ�GE ����o��6�!E EN0�A�_��v{�y|��q����D4^a"A4�6^�2��F
rȟ*��Z�R!튉#]���(`m@t�6!YH���yY ��3�&��gH�8�*��#���CsU"�)�J��E�+-��N#X�Fl�2�72�t!�F�\���R#J(���/(��G�����{lc��A
~�;:�����8K�u�P��"��`�K�AsE�k��P�S��sɶEFE�t��$��ɏ�ʵ&���FQ2b��_f=Jc/����/d��H�16#�'����W[�(����-Hj _P��"�s[�}'��)왔��E���ƌZ9]���f���`a��20/������ �����tБ�@�w��oJ%g�_�܃:��hl� ���c�g����D�`=F&�S��G��7q^Oy�C�l�~�.5�sy�ɢ�:"*L���U�"Bx�^"m�� l����<;���
�"W���˴�hv#Rr�	I9��;y���@�T���Ci��t�C
���Rah1(AC��W%Ԙ�&" hm��,��	���p1^���vưcЖ�K�*��ȸ+ޗ.!���(U��kC�IB9)j��9W`Q׽L�-�g��K�A��U�H;�q
���q(�1�-��?"d�#I9���n bl`؆=7�����J/՟/�rY�p���#�+�RKD#`��샠cI��^>@< sJ�p��/�H*��hhm^��Ǩ���#@��.�	 8APR0�����#�	o���4XdP- c��D����̓��l.�+$eMH5��v�D�1�@h@S�1�@���vG����D���X���i80�\�� &��t�{�j��?>���� LI��I��| ��Q��%��.7��;�ܩ�)d���e �P:9�	 �M���Ӂ�KKB��.�{ɫs��rT�H�_ʇ��IK'����`�%:��Ϊ��d��)��Fsf��ֲ͎h7����,�H4w�4����`L:�L��a�!#X�b��erP�.sy��fcA�6����9��3��$#��7~�1?���)���